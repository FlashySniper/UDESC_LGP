<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-12.991,-25.1033,145.053,-105.903</PageViewport>
<gate>
<ID>2</ID>
<type>AA_LABEL</type>
<position>5,-7</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>4</ID>
<type>AA_LABEL</type>
<position>9,-7</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>5</ID>
<type>AA_LABEL</type>
<position>12.5,-7</position>
<gparam>LABEL_TEXT S</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>7</ID>
<type>AA_LABEL</type>
<position>5,-10.5</position>
<gparam>LABEL_TEXT 0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>8</ID>
<type>AA_LABEL</type>
<position>5,-13.5</position>
<gparam>LABEL_TEXT 0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>9</ID>
<type>AA_LABEL</type>
<position>5,-16.5</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>10</ID>
<type>AA_LABEL</type>
<position>5,-19.5</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>11</ID>
<type>AA_LABEL</type>
<position>9,-19.5</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>15</ID>
<type>AI_XOR2</type>
<position>41.5,-14</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>17</ID>
<type>AA_TOGGLE</type>
<position>29.5,-12.5</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>19</ID>
<type>AA_TOGGLE</type>
<position>29.5,-15.5</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>22</ID>
<type>AA_LABEL</type>
<position>9,-13.5</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>23</ID>
<type>AA_LABEL</type>
<position>9,-16.5</position>
<gparam>LABEL_TEXT 0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>24</ID>
<type>AA_LABEL</type>
<position>9,-10.5</position>
<gparam>LABEL_TEXT 0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>25</ID>
<type>AA_LABEL</type>
<position>12.5,-19.5</position>
<gparam>LABEL_TEXT 0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>26</ID>
<type>AA_LABEL</type>
<position>12.5,-10.5</position>
<gparam>LABEL_TEXT 0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>28</ID>
<type>AA_LABEL</type>
<position>12.5,-13.5</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>29</ID>
<type>AA_LABEL</type>
<position>12.5,-16.5</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>31</ID>
<type>AI_XOR2</type>
<position>54.5,-15</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>4 </input>
<output>
<ID>OUT</ID>5 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>33</ID>
<type>AA_TOGGLE</type>
<position>29.5,-18.5</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>34</ID>
<type>AA_LABEL</type>
<position>26.5,-12</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>36</ID>
<type>AA_LABEL</type>
<position>26.5,-15</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>37</ID>
<type>AA_LABEL</type>
<position>26.5,-18</position>
<gparam>LABEL_TEXT C</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>39</ID>
<type>GA_LED</type>
<position>62,-15</position>
<input>
<ID>N_in0</ID>5 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>40</ID>
<type>AA_LABEL</type>
<position>62,-11.5</position>
<gparam>LABEL_TEXT S</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>44</ID>
<type>AA_AND2</type>
<position>37.5,-27</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>46</ID>
<type>AE_OR2</type>
<position>57,-29</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>7 </input>
<output>
<ID>OUT</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>48</ID>
<type>AA_AND2</type>
<position>50.5,-23.5</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>3 </input>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>50</ID>
<type>GA_LED</type>
<position>66,-29</position>
<input>
<ID>N_in0</ID>9 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>52</ID>
<type>AA_LABEL</type>
<position>71,-28.5</position>
<gparam>LABEL_TEXT Cout</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>56</ID>
<type>AA_TOGGLE</type>
<position>5,-37</position>
<output>
<ID>OUT_0</ID>44 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>57</ID>
<type>AA_TOGGLE</type>
<position>8,-37</position>
<output>
<ID>OUT_0</ID>38 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>58</ID>
<type>AA_TOGGLE</type>
<position>11,-37</position>
<output>
<ID>OUT_0</ID>30 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>59</ID>
<type>AA_TOGGLE</type>
<position>14,-37</position>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>60</ID>
<type>AA_TOGGLE</type>
<position>22.5,-37</position>
<output>
<ID>OUT_0</ID>43 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>61</ID>
<type>AA_TOGGLE</type>
<position>25,-37</position>
<output>
<ID>OUT_0</ID>37 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>62</ID>
<type>AA_TOGGLE</type>
<position>28,-37</position>
<output>
<ID>OUT_0</ID>29 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>63</ID>
<type>AA_TOGGLE</type>
<position>31.5,-37</position>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>64</ID>
<type>AA_LABEL</type>
<position>5,-34.5</position>
<gparam>LABEL_TEXT A3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>65</ID>
<type>AA_LABEL</type>
<position>8,-34.5</position>
<gparam>LABEL_TEXT A2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>66</ID>
<type>AA_LABEL</type>
<position>11,-34.5</position>
<gparam>LABEL_TEXT A1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>67</ID>
<type>AA_LABEL</type>
<position>14,-34.5</position>
<gparam>LABEL_TEXT A0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>68</ID>
<type>AA_LABEL</type>
<position>31,-34.5</position>
<gparam>LABEL_TEXT B0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>69</ID>
<type>AA_LABEL</type>
<position>28,-34.5</position>
<gparam>LABEL_TEXT B1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>70</ID>
<type>AA_LABEL</type>
<position>25,-34.5</position>
<gparam>LABEL_TEXT B2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>71</ID>
<type>AA_LABEL</type>
<position>22,-34.5</position>
<gparam>LABEL_TEXT B3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>73</ID>
<type>AI_XOR2</type>
<position>41,-46</position>
<input>
<ID>IN_0</ID>10 </input>
<input>
<ID>IN_1</ID>11 </input>
<output>
<ID>OUT</ID>25 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>81</ID>
<type>GA_LED</type>
<position>68,-46.5</position>
<input>
<ID>N_in0</ID>26 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>82</ID>
<type>AA_LABEL</type>
<position>68,-44.5</position>
<gparam>LABEL_TEXT S0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>90</ID>
<type>GA_LED</type>
<position>75.5,-62.5</position>
<input>
<ID>N_in0</ID>33 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>91</ID>
<type>AA_LABEL</type>
<position>75.5,-59.5</position>
<gparam>LABEL_TEXT S1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>99</ID>
<type>AA_TOGGLE</type>
<position>36,-40</position>
<output>
<ID>OUT_0</ID>24 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>101</ID>
<type>AI_XOR2</type>
<position>53,-47.5</position>
<input>
<ID>IN_0</ID>25 </input>
<input>
<ID>IN_1</ID>24 </input>
<output>
<ID>OUT</ID>26 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>103</ID>
<type>AA_AND2</type>
<position>47,-55.5</position>
<input>
<ID>IN_0</ID>25 </input>
<input>
<ID>IN_1</ID>24 </input>
<output>
<ID>OUT</ID>27 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>104</ID>
<type>AA_LABEL</type>
<position>36,-38</position>
<gparam>LABEL_TEXT C</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>106</ID>
<type>AA_AND2</type>
<position>47,-61.5</position>
<input>
<ID>IN_0</ID>10 </input>
<input>
<ID>IN_1</ID>11 </input>
<output>
<ID>OUT</ID>28 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>108</ID>
<type>AE_OR2</type>
<position>57.5,-59</position>
<input>
<ID>IN_0</ID>27 </input>
<input>
<ID>IN_1</ID>28 </input>
<output>
<ID>OUT</ID>31 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>110</ID>
<type>AI_XOR2</type>
<position>58,-69</position>
<input>
<ID>IN_0</ID>29 </input>
<input>
<ID>IN_1</ID>30 </input>
<output>
<ID>OUT</ID>32 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>112</ID>
<type>AI_XOR2</type>
<position>68,-62.5</position>
<input>
<ID>IN_0</ID>31 </input>
<input>
<ID>IN_1</ID>32 </input>
<output>
<ID>OUT</ID>33 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>113</ID>
<type>AA_LABEL</type>
<position>57,-55.5</position>
<gparam>LABEL_TEXT C</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>115</ID>
<type>AA_AND2</type>
<position>66.5,-77.5</position>
<input>
<ID>IN_0</ID>31 </input>
<input>
<ID>IN_1</ID>32 </input>
<output>
<ID>OUT</ID>34 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>117</ID>
<type>AA_AND2</type>
<position>67,-84</position>
<input>
<ID>IN_0</ID>29 </input>
<input>
<ID>IN_1</ID>30 </input>
<output>
<ID>OUT</ID>35 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>119</ID>
<type>AE_OR2</type>
<position>75.5,-80.5</position>
<input>
<ID>IN_0</ID>34 </input>
<input>
<ID>IN_1</ID>35 </input>
<output>
<ID>OUT</ID>36 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>120</ID>
<type>AA_LABEL</type>
<position>75,-76.5</position>
<gparam>LABEL_TEXT C</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>122</ID>
<type>AI_XOR2</type>
<position>88.5,-81.5</position>
<input>
<ID>IN_0</ID>36 </input>
<input>
<ID>IN_1</ID>39 </input>
<output>
<ID>OUT</ID>40 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>124</ID>
<type>AI_XOR2</type>
<position>82,-89</position>
<input>
<ID>IN_0</ID>37 </input>
<input>
<ID>IN_1</ID>38 </input>
<output>
<ID>OUT</ID>39 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>125</ID>
<type>GA_LED</type>
<position>96,-82</position>
<input>
<ID>N_in0</ID>40 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>126</ID>
<type>AA_LABEL</type>
<position>96,-79.5</position>
<gparam>LABEL_TEXT S2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>128</ID>
<type>AA_AND2</type>
<position>90,-95.5</position>
<input>
<ID>IN_0</ID>39 </input>
<input>
<ID>IN_1</ID>36 </input>
<output>
<ID>OUT</ID>41 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>130</ID>
<type>AA_AND2</type>
<position>90,-101.5</position>
<input>
<ID>IN_0</ID>37 </input>
<input>
<ID>IN_1</ID>38 </input>
<output>
<ID>OUT</ID>42 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>132</ID>
<type>AE_OR2</type>
<position>99,-98.5</position>
<input>
<ID>IN_0</ID>41 </input>
<input>
<ID>IN_1</ID>42 </input>
<output>
<ID>OUT</ID>45 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>133</ID>
<type>AA_LABEL</type>
<position>98.5,-95</position>
<gparam>LABEL_TEXT C</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>135</ID>
<type>AA_FULLADDER_1BIT</type>
<position>112.5,-95</position>
<input>
<ID>IN_0</ID>43 </input>
<input>
<ID>IN_B_0</ID>44 </input>
<output>
<ID>OUT_0</ID>46 </output>
<input>
<ID>carry_in</ID>45 </input>
<output>
<ID>carry_out</ID>47 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>136</ID>
<type>GA_LED</type>
<position>120,-98.5</position>
<input>
<ID>N_in0</ID>46 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>137</ID>
<type>AA_LABEL</type>
<position>120,-96</position>
<gparam>LABEL_TEXT S3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>138</ID>
<type>GA_LED</type>
<position>106,-95</position>
<input>
<ID>N_in1</ID>47 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>139</ID>
<type>AA_LABEL</type>
<position>106,-92.5</position>
<gparam>LABEL_TEXT S4</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31.5,-12.5,34,-12.5</points>
<connection>
<GID>17</GID>
<name>OUT_0</name></connection>
<intersection>34 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>34,-26,34,-12.5</points>
<intersection>-26 10</intersection>
<intersection>-13 8</intersection>
<intersection>-12.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>34,-13,38.5,-13</points>
<connection>
<GID>15</GID>
<name>IN_0</name></connection>
<intersection>34 6</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>34,-26,34.5,-26</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<intersection>34 6</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31.5,-15.5,33,-15.5</points>
<connection>
<GID>19</GID>
<name>OUT_0</name></connection>
<intersection>33 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>33,-28,33,-15</points>
<intersection>-28 9</intersection>
<intersection>-15.5 1</intersection>
<intersection>-15 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>33,-15,38.5,-15</points>
<connection>
<GID>15</GID>
<name>IN_1</name></connection>
<intersection>33 4</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>33,-28,34.5,-28</points>
<connection>
<GID>44</GID>
<name>IN_1</name></connection>
<intersection>33 4</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>44.5,-24.5,44.5,-14</points>
<intersection>-24.5 8</intersection>
<intersection>-14 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>44.5,-14,51.5,-14</points>
<connection>
<GID>15</GID>
<name>OUT</name></connection>
<connection>
<GID>31</GID>
<name>IN_0</name></connection>
<intersection>44.5 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>44.5,-24.5,47.5,-24.5</points>
<connection>
<GID>48</GID>
<name>IN_1</name></connection>
<intersection>44.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46,-22.5,46,-16</points>
<intersection>-22.5 4</intersection>
<intersection>-18.5 2</intersection>
<intersection>-16 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46,-16,51.5,-16</points>
<connection>
<GID>31</GID>
<name>IN_1</name></connection>
<intersection>46 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>31.5,-18.5,46,-18.5</points>
<connection>
<GID>33</GID>
<name>OUT_0</name></connection>
<intersection>46 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>46,-22.5,47.5,-22.5</points>
<connection>
<GID>48</GID>
<name>IN_0</name></connection>
<intersection>46 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57.5,-15,61,-15</points>
<connection>
<GID>39</GID>
<name>N_in0</name></connection>
<connection>
<GID>31</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40.5,-30,54,-30</points>
<connection>
<GID>46</GID>
<name>IN_1</name></connection>
<intersection>40.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>40.5,-30,40.5,-27</points>
<connection>
<GID>44</GID>
<name>OUT</name></connection>
<intersection>-30 1</intersection></vsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53.5,-28,53.5,-23.5</points>
<connection>
<GID>48</GID>
<name>OUT</name></connection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>53.5,-28,54,-28</points>
<connection>
<GID>46</GID>
<name>IN_0</name></connection>
<intersection>53.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>60,-29,65,-29</points>
<connection>
<GID>50</GID>
<name>N_in0</name></connection>
<connection>
<GID>46</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31.5,-60.5,31.5,-39</points>
<connection>
<GID>63</GID>
<name>OUT_0</name></connection>
<intersection>-60.5 5</intersection>
<intersection>-45 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31.5,-45,38,-45</points>
<connection>
<GID>73</GID>
<name>IN_0</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>31.5,-60.5,44,-60.5</points>
<connection>
<GID>106</GID>
<name>IN_0</name></connection>
<intersection>31.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14,-62.5,14,-39</points>
<connection>
<GID>59</GID>
<name>OUT_0</name></connection>
<intersection>-62.5 5</intersection>
<intersection>-47 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>14,-47,38,-47</points>
<connection>
<GID>73</GID>
<name>IN_1</name></connection>
<intersection>14 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>14,-62.5,44,-62.5</points>
<connection>
<GID>106</GID>
<name>IN_1</name></connection>
<intersection>14 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,-56.5,36,-42</points>
<connection>
<GID>99</GID>
<name>OUT_0</name></connection>
<intersection>-56.5 3</intersection>
<intersection>-48.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36,-48.5,50,-48.5</points>
<connection>
<GID>101</GID>
<name>IN_1</name></connection>
<intersection>36 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>36,-56.5,44,-56.5</points>
<connection>
<GID>103</GID>
<name>IN_1</name></connection>
<intersection>36 0</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47,-46.5,47,-46</points>
<intersection>-46.5 1</intersection>
<intersection>-46 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,-46.5,50,-46.5</points>
<connection>
<GID>101</GID>
<name>IN_0</name></connection>
<intersection>47 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>44,-46,47,-46</points>
<connection>
<GID>73</GID>
<name>OUT</name></connection>
<intersection>44 3</intersection>
<intersection>47 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>44,-54.5,44,-46</points>
<connection>
<GID>103</GID>
<name>IN_0</name></connection>
<intersection>-46 2</intersection></vsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61.5,-47.5,61.5,-46.5</points>
<intersection>-47.5 2</intersection>
<intersection>-46.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>61.5,-46.5,67,-46.5</points>
<connection>
<GID>81</GID>
<name>N_in0</name></connection>
<intersection>61.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56,-47.5,61.5,-47.5</points>
<connection>
<GID>101</GID>
<name>OUT</name></connection>
<intersection>61.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52,-58,52,-55.5</points>
<intersection>-58 1</intersection>
<intersection>-55.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>52,-58,54.5,-58</points>
<connection>
<GID>108</GID>
<name>IN_0</name></connection>
<intersection>52 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>50,-55.5,52,-55.5</points>
<connection>
<GID>103</GID>
<name>OUT</name></connection>
<intersection>52 0</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52,-61.5,52,-60</points>
<intersection>-61.5 2</intersection>
<intersection>-60 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>52,-60,54.5,-60</points>
<connection>
<GID>108</GID>
<name>IN_1</name></connection>
<intersection>52 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>50,-61.5,52,-61.5</points>
<connection>
<GID>106</GID>
<name>OUT</name></connection>
<intersection>52 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,-68,28,-39</points>
<connection>
<GID>62</GID>
<name>OUT_0</name></connection>
<intersection>-68 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28,-68,55,-68</points>
<connection>
<GID>110</GID>
<name>IN_0</name></connection>
<intersection>28 0</intersection>
<intersection>52.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>52.5,-83,52.5,-68</points>
<intersection>-83 3</intersection>
<intersection>-68 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>52.5,-83,64,-83</points>
<connection>
<GID>117</GID>
<name>IN_0</name></connection>
<intersection>52.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11,-70,11,-39</points>
<connection>
<GID>58</GID>
<name>OUT_0</name></connection>
<intersection>-70 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>11,-70,55,-70</points>
<connection>
<GID>110</GID>
<name>IN_1</name></connection>
<intersection>11 0</intersection>
<intersection>49 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>49,-85,49,-70</points>
<intersection>-85 3</intersection>
<intersection>-70 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>49,-85,64,-85</points>
<connection>
<GID>117</GID>
<name>IN_1</name></connection>
<intersection>49 2</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61.5,-76.5,61.5,-59</points>
<intersection>-76.5 4</intersection>
<intersection>-61.5 3</intersection>
<intersection>-59 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>60.5,-59,61.5,-59</points>
<connection>
<GID>108</GID>
<name>OUT</name></connection>
<intersection>61.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>61.5,-61.5,65,-61.5</points>
<connection>
<GID>112</GID>
<name>IN_0</name></connection>
<intersection>61.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>61.5,-76.5,63.5,-76.5</points>
<connection>
<GID>115</GID>
<name>IN_0</name></connection>
<intersection>61.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62.5,-78.5,62.5,-63.5</points>
<intersection>-78.5 5</intersection>
<intersection>-69 2</intersection>
<intersection>-63.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>61,-69,62.5,-69</points>
<connection>
<GID>110</GID>
<name>OUT</name></connection>
<intersection>62.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>62.5,-63.5,65,-63.5</points>
<connection>
<GID>112</GID>
<name>IN_1</name></connection>
<intersection>62.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>62.5,-78.5,63.5,-78.5</points>
<connection>
<GID>115</GID>
<name>IN_1</name></connection>
<intersection>62.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71,-62.5,74.5,-62.5</points>
<connection>
<GID>90</GID>
<name>N_in0</name></connection>
<connection>
<GID>112</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>71,-79.5,71,-77.5</points>
<intersection>-79.5 1</intersection>
<intersection>-77.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>71,-79.5,72.5,-79.5</points>
<connection>
<GID>119</GID>
<name>IN_0</name></connection>
<intersection>71 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>69.5,-77.5,71,-77.5</points>
<connection>
<GID>115</GID>
<name>OUT</name></connection>
<intersection>71 0</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>71,-84,71,-81.5</points>
<intersection>-84 2</intersection>
<intersection>-81.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>71,-81.5,72.5,-81.5</points>
<connection>
<GID>119</GID>
<name>IN_1</name></connection>
<intersection>71 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>70,-84,71,-84</points>
<connection>
<GID>117</GID>
<name>OUT</name></connection>
<intersection>71 0</intersection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78.5,-80.5,85.5,-80.5</points>
<connection>
<GID>119</GID>
<name>OUT</name></connection>
<connection>
<GID>122</GID>
<name>IN_0</name></connection>
<intersection>84.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>84.5,-96.5,84.5,-80.5</points>
<intersection>-96.5 7</intersection>
<intersection>-80.5 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>84.5,-96.5,87,-96.5</points>
<connection>
<GID>128</GID>
<name>IN_1</name></connection>
<intersection>84.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,-88,25,-39</points>
<connection>
<GID>61</GID>
<name>OUT_0</name></connection>
<intersection>-88 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25,-88,79,-88</points>
<connection>
<GID>124</GID>
<name>IN_0</name></connection>
<intersection>25 0</intersection>
<intersection>73 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>73,-100.5,73,-88</points>
<intersection>-100.5 3</intersection>
<intersection>-88 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>73,-100.5,87,-100.5</points>
<connection>
<GID>130</GID>
<name>IN_0</name></connection>
<intersection>73 2</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8,-90,8,-39</points>
<connection>
<GID>57</GID>
<name>OUT_0</name></connection>
<intersection>-90 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>8,-90,79,-90</points>
<connection>
<GID>124</GID>
<name>IN_1</name></connection>
<intersection>8 0</intersection>
<intersection>71.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>71.5,-102.5,71.5,-90</points>
<intersection>-102.5 3</intersection>
<intersection>-90 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>71.5,-102.5,87,-102.5</points>
<connection>
<GID>130</GID>
<name>IN_1</name></connection>
<intersection>71.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85,-94.5,85,-82.5</points>
<connection>
<GID>124</GID>
<name>OUT</name></connection>
<intersection>-94.5 2</intersection>
<intersection>-82.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>85,-82.5,85.5,-82.5</points>
<connection>
<GID>122</GID>
<name>IN_1</name></connection>
<intersection>85 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>85,-94.5,87,-94.5</points>
<connection>
<GID>128</GID>
<name>IN_0</name></connection>
<intersection>85 0</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>93,-82,93,-81.5</points>
<intersection>-82 1</intersection>
<intersection>-81.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>93,-82,95,-82</points>
<connection>
<GID>125</GID>
<name>N_in0</name></connection>
<intersection>93 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>91.5,-81.5,93,-81.5</points>
<connection>
<GID>122</GID>
<name>OUT</name></connection>
<intersection>93 0</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>94.5,-97.5,94.5,-95.5</points>
<intersection>-97.5 1</intersection>
<intersection>-95.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>94.5,-97.5,96,-97.5</points>
<connection>
<GID>132</GID>
<name>IN_0</name></connection>
<intersection>94.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>93,-95.5,94.5,-95.5</points>
<connection>
<GID>128</GID>
<name>OUT</name></connection>
<intersection>94.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>94.5,-101.5,94.5,-99.5</points>
<intersection>-101.5 2</intersection>
<intersection>-99.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>94.5,-99.5,96,-99.5</points>
<connection>
<GID>132</GID>
<name>IN_1</name></connection>
<intersection>94.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>93,-101.5,94.5,-101.5</points>
<connection>
<GID>130</GID>
<name>OUT</name></connection>
<intersection>94.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>113.5,-92,113.5,-68</points>
<connection>
<GID>135</GID>
<name>IN_0</name></connection>
<intersection>-68 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>22.5,-68,22.5,-39</points>
<connection>
<GID>60</GID>
<name>OUT_0</name></connection>
<intersection>-68 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>22.5,-68,113.5,-68</points>
<intersection>22.5 1</intersection>
<intersection>113.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111.5,-92,111.5,-68</points>
<connection>
<GID>135</GID>
<name>IN_B_0</name></connection>
<intersection>-68 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>5,-68,5,-39</points>
<connection>
<GID>56</GID>
<name>OUT_0</name></connection>
<intersection>-68 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>5,-68,111.5,-68</points>
<intersection>5 1</intersection>
<intersection>111.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>102,-101,116.5,-101</points>
<intersection>102 3</intersection>
<intersection>116.5 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>102,-101,102,-98.5</points>
<connection>
<GID>132</GID>
<name>OUT</name></connection>
<intersection>-101 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>116.5,-101,116.5,-95</points>
<connection>
<GID>135</GID>
<name>carry_in</name></connection>
<intersection>-101 1</intersection></vsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>112.5,-98.5,112.5,-98</points>
<connection>
<GID>135</GID>
<name>OUT_0</name></connection>
<intersection>-98.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>112.5,-98.5,119,-98.5</points>
<connection>
<GID>136</GID>
<name>N_in0</name></connection>
<intersection>112.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>107,-95,108.5,-95</points>
<connection>
<GID>138</GID>
<name>N_in1</name></connection>
<connection>
<GID>135</GID>
<name>carry_out</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,177.8,-90.9</PageViewport></page 1>
<page 2>
<PageViewport>0,0,177.8,-90.9</PageViewport></page 2>
<page 3>
<PageViewport>0,0,177.8,-90.9</PageViewport></page 3>
<page 4>
<PageViewport>0,0,177.8,-90.9</PageViewport></page 4>
<page 5>
<PageViewport>0,0,177.8,-90.9</PageViewport></page 5>
<page 6>
<PageViewport>0,0,177.8,-90.9</PageViewport></page 6>
<page 7>
<PageViewport>0,0,177.8,-90.9</PageViewport></page 7>
<page 8>
<PageViewport>0,0,177.8,-90.9</PageViewport></page 8>
<page 9>
<PageViewport>0,0,177.8,-90.9</PageViewport></page 9></circuit>